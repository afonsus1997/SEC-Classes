

module push_button_driver(
    input sel,
    input [3:0] sw_in,
    output [3:0], sw_out
);

endmodule // push_button_driver