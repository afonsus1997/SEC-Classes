

module sequencer_loop_ctl(
    input [7:0] freq,
    input [7:0] kbd_in.
    input sel_loop,
    input sel_snd,
    output snd_out,
    output reg [7:0] led_out
);




endmodule // sequencerloopctl
