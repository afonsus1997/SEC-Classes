

module led_driver(
    input [7:0] data_in,
    output [7:0] led_out
);

endmodule // led_driver