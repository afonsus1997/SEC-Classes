

module switch_driver(
    input sel,
    input [7:0] kbd_in,
    output [7:0] kbd_out
    output [7:0] led_out
);

endmodule // switch_driver